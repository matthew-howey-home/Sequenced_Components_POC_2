
module Internal_Oscillator (
	clkout,
	oscena);	

	output		clkout;
	input		oscena;
endmodule
